CDLv2�H�\                                                                                                                   				    		                                                                                                     	                     	                                                                                                                                                                                                                                                                                                                 	                                         	                                                                                                                                           	                                                                           		            	                                				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    							      		         		                      	     	                                                                                                                                                                                                                                                                                                     				                                                                                                                                                                                                                                                  	                                      		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        	                                                                                                                                                                                                                                                                                                                                                                                                                                                            	                                                                    			                  	             				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    	  		                                                                                                                                                                                                                                                                                               	   	                                                                                                                                     	                                                                                                                                        	                                                                               			                                                                        	                                                                                                                                   	                                         	                                                                                                                                                       	                                                                                                                                                                                                                                                                                                                                                           	                                                                                                                                                                                                                                                                                                                                                                             	       	         	            			                  	                           		                         	                              	                                                            	                                                   					                                          	                                                                              	                                                                                                                                                                                                                                                    	           	                                                                                                                                                                                         	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      	                                                                                                                                                                                                                                                                      	                                                          	                                                                         	           		                                                                           	                                                                                                                                                                                                                                                            			                                                                                                                                                                                                                                                                                		                   	 	                                                                                            	           	 		     	        	                                                                                                                                                                                                                       		                                                                           			                                     			               	   		                                    	                     				                                                                                                                                                                                                                                                                                                                                                                                                         		                                                                                                                                             	               	                                                                                                                                                                                                                                                                                                                                                 	                                                                                                                                                                                                                                                                                                                                                                                                   		          		                 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           	                                                                                     			                                				          							          	 					  	      					   		                                    	                                                                                                                                                                                                                                                                               	                                                                                                                                                           	                                 	                                                                                           			      	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      